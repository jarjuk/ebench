[HEAD]:115
VPP:2.400000
OFFSET:0.000000
CHANNEL:1
RATEPOS:0.000031
RATENEG:0.000031
MAX:32767.000000
MIN:-32767.000000
[DATA]:0
